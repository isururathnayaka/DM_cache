// Content          : Cache controller
// Author           : Isuru Rathnayaka
// Last Modified    : 2019.09.13

import memory_sub_system_config::*;

module cache_controller();


endmodule

